module Random(output reg [1:0] num1, num2, input [4:0] seqNo, input [5:0] idx1, idx2);



reg seq[19:0][49:0][1:0];




always@(*)
begin
num1 = {seq[seqNo][idx1][1],seq[seqNo][idx1][0]};
num2 = {seq[seqNo][idx2][1],seq[seqNo][idx2][0]};
end


initial
begin
seq[0][0][0] = 1'b0;
seq[0][0][1] = 1'b0;
seq[0][1][0] = 1'b1;
seq[0][1][1] = 1'b1;
seq[0][2][0] = 1'b1;
seq[0][2][1] = 1'b0;
seq[0][3][0] = 1'b1;
seq[0][3][1] = 1'b1;
seq[0][4][0] = 1'b0;
seq[0][4][1] = 1'b0;
seq[0][5][0] = 1'b0;
seq[0][5][1] = 1'b1;
seq[0][6][0] = 1'b1;
seq[0][6][1] = 1'b1;
seq[0][7][0] = 1'b0;
seq[0][7][1] = 1'b0;
seq[0][8][0] = 1'b1;
seq[0][8][1] = 1'b0;
seq[0][9][0] = 1'b1;
seq[0][9][1] = 1'b1;
seq[0][10][0] = 1'b1;
seq[0][10][1] = 1'b0;
seq[0][11][0] = 1'b0;
seq[0][11][1] = 1'b1;
seq[0][12][0] = 1'b1;
seq[0][12][1] = 1'b0;
seq[0][13][0] = 1'b0;
seq[0][13][1] = 1'b1;
seq[0][14][0] = 1'b0;
seq[0][14][1] = 1'b1;
seq[0][15][0] = 1'b0;
seq[0][15][1] = 1'b1;
seq[0][16][0] = 1'b1;
seq[0][16][1] = 1'b1;
seq[0][17][0] = 1'b0;
seq[0][17][1] = 1'b1;
seq[0][18][0] = 1'b1;
seq[0][18][1] = 1'b0;
seq[0][19][0] = 1'b1;
seq[0][19][1] = 1'b0;
seq[0][20][0] = 1'b0;
seq[0][20][1] = 1'b0;
seq[0][21][0] = 1'b0;
seq[0][21][1] = 1'b0;
seq[0][22][0] = 1'b1;
seq[0][22][1] = 1'b1;
seq[0][23][0] = 1'b0;
seq[0][23][1] = 1'b0;
seq[0][24][0] = 1'b0;
seq[0][24][1] = 1'b1;
seq[0][25][0] = 1'b1;
seq[0][25][1] = 1'b0;
seq[0][26][0] = 1'b0;
seq[0][26][1] = 1'b1;
seq[0][27][0] = 1'b1;
seq[0][27][1] = 1'b0;
seq[0][28][0] = 1'b0;
seq[0][28][1] = 1'b0;
seq[0][29][0] = 1'b0;
seq[0][29][1] = 1'b1;
seq[0][30][0] = 1'b1;
seq[0][30][1] = 1'b0;
seq[0][31][0] = 1'b0;
seq[0][31][1] = 1'b0;
seq[0][32][0] = 1'b1;
seq[0][32][1] = 1'b0;
seq[0][33][0] = 1'b0;
seq[0][33][1] = 1'b0;
seq[0][34][0] = 1'b0;
seq[0][34][1] = 1'b1;
seq[0][35][0] = 1'b1;
seq[0][35][1] = 1'b1;
seq[0][36][0] = 1'b0;
seq[0][36][1] = 1'b1;
seq[0][37][0] = 1'b1;
seq[0][37][1] = 1'b0;
seq[0][38][0] = 1'b1;
seq[0][38][1] = 1'b0;
seq[0][39][0] = 1'b1;
seq[0][39][1] = 1'b0;
seq[0][40][0] = 1'b1;
seq[0][40][1] = 1'b0;
seq[0][41][0] = 1'b0;
seq[0][41][1] = 1'b1;
seq[0][42][0] = 1'b0;
seq[0][42][1] = 1'b1;
seq[0][43][0] = 1'b0;
seq[0][43][1] = 1'b0;
seq[0][44][0] = 1'b1;
seq[0][44][1] = 1'b1;
seq[0][45][0] = 1'b0;
seq[0][45][1] = 1'b0;
seq[0][46][0] = 1'b1;
seq[0][46][1] = 1'b0;
seq[0][47][0] = 1'b0;
seq[0][47][1] = 1'b0;
seq[0][48][0] = 1'b0;
seq[0][48][1] = 1'b1;
seq[0][49][0] = 1'b0;
seq[0][49][1] = 1'b0;
seq[1][0][0] = 1'b0;
seq[1][0][1] = 1'b0;
seq[1][1][0] = 1'b0;
seq[1][1][1] = 1'b1;
seq[1][2][0] = 1'b0;
seq[1][2][1] = 1'b1;
seq[1][3][0] = 1'b1;
seq[1][3][1] = 1'b1;
seq[1][4][0] = 1'b0;
seq[1][4][1] = 1'b0;
seq[1][5][0] = 1'b1;
seq[1][5][1] = 1'b1;
seq[1][6][0] = 1'b1;
seq[1][6][1] = 1'b0;
seq[1][7][0] = 1'b1;
seq[1][7][1] = 1'b1;
seq[1][8][0] = 1'b1;
seq[1][8][1] = 1'b0;
seq[1][9][0] = 1'b0;
seq[1][9][1] = 1'b0;
seq[1][10][0] = 1'b0;
seq[1][10][1] = 1'b0;
seq[1][11][0] = 1'b1;
seq[1][11][1] = 1'b1;
seq[1][12][0] = 1'b0;
seq[1][12][1] = 1'b0;
seq[1][13][0] = 1'b0;
seq[1][13][1] = 1'b0;
seq[1][14][0] = 1'b1;
seq[1][14][1] = 1'b1;
seq[1][15][0] = 1'b0;
seq[1][15][1] = 1'b0;
seq[1][16][0] = 1'b0;
seq[1][16][1] = 1'b0;
seq[1][17][0] = 1'b1;
seq[1][17][1] = 1'b1;
seq[1][18][0] = 1'b1;
seq[1][18][1] = 1'b1;
seq[1][19][0] = 1'b1;
seq[1][19][1] = 1'b1;
seq[1][20][0] = 1'b1;
seq[1][20][1] = 1'b0;
seq[1][21][0] = 1'b0;
seq[1][21][1] = 1'b1;
seq[1][22][0] = 1'b0;
seq[1][22][1] = 1'b0;
seq[1][23][0] = 1'b1;
seq[1][23][1] = 1'b1;
seq[1][24][0] = 1'b1;
seq[1][24][1] = 1'b1;
seq[1][25][0] = 1'b0;
seq[1][25][1] = 1'b0;
seq[1][26][0] = 1'b1;
seq[1][26][1] = 1'b1;
seq[1][27][0] = 1'b0;
seq[1][27][1] = 1'b1;
seq[1][28][0] = 1'b1;
seq[1][28][1] = 1'b0;
seq[1][29][0] = 1'b0;
seq[1][29][1] = 1'b1;
seq[1][30][0] = 1'b0;
seq[1][30][1] = 1'b1;
seq[1][31][0] = 1'b1;
seq[1][31][1] = 1'b1;
seq[1][32][0] = 1'b0;
seq[1][32][1] = 1'b1;
seq[1][33][0] = 1'b1;
seq[1][33][1] = 1'b0;
seq[1][34][0] = 1'b1;
seq[1][34][1] = 1'b1;
seq[1][35][0] = 1'b0;
seq[1][35][1] = 1'b1;
seq[1][36][0] = 1'b1;
seq[1][36][1] = 1'b1;
seq[1][37][0] = 1'b0;
seq[1][37][1] = 1'b0;
seq[1][38][0] = 1'b0;
seq[1][38][1] = 1'b1;
seq[1][39][0] = 1'b0;
seq[1][39][1] = 1'b0;
seq[1][40][0] = 1'b0;
seq[1][40][1] = 1'b0;
seq[1][41][0] = 1'b1;
seq[1][41][1] = 1'b1;
seq[1][42][0] = 1'b1;
seq[1][42][1] = 1'b0;
seq[1][43][0] = 1'b0;
seq[1][43][1] = 1'b0;
seq[1][44][0] = 1'b0;
seq[1][44][1] = 1'b0;
seq[1][45][0] = 1'b1;
seq[1][45][1] = 1'b0;
seq[1][46][0] = 1'b0;
seq[1][46][1] = 1'b0;
seq[1][47][0] = 1'b0;
seq[1][47][1] = 1'b0;
seq[1][48][0] = 1'b1;
seq[1][48][1] = 1'b1;
seq[1][49][0] = 1'b1;
seq[1][49][1] = 1'b1;
seq[2][0][0] = 1'b0;
seq[2][0][1] = 1'b0;
seq[2][1][0] = 1'b0;
seq[2][1][1] = 1'b0;
seq[2][2][0] = 1'b1;
seq[2][2][1] = 1'b0;
seq[2][3][0] = 1'b1;
seq[2][3][1] = 1'b0;
seq[2][4][0] = 1'b0;
seq[2][4][1] = 1'b0;
seq[2][5][0] = 1'b0;
seq[2][5][1] = 1'b1;
seq[2][6][0] = 1'b1;
seq[2][6][1] = 1'b0;
seq[2][7][0] = 1'b0;
seq[2][7][1] = 1'b0;
seq[2][8][0] = 1'b0;
seq[2][8][1] = 1'b1;
seq[2][9][0] = 1'b1;
seq[2][9][1] = 1'b1;
seq[2][10][0] = 1'b1;
seq[2][10][1] = 1'b1;
seq[2][11][0] = 1'b1;
seq[2][11][1] = 1'b1;
seq[2][12][0] = 1'b0;
seq[2][12][1] = 1'b0;
seq[2][13][0] = 1'b1;
seq[2][13][1] = 1'b0;
seq[2][14][0] = 1'b0;
seq[2][14][1] = 1'b0;
seq[2][15][0] = 1'b0;
seq[2][15][1] = 1'b0;
seq[2][16][0] = 1'b0;
seq[2][16][1] = 1'b0;
seq[2][17][0] = 1'b1;
seq[2][17][1] = 1'b0;
seq[2][18][0] = 1'b0;
seq[2][18][1] = 1'b0;
seq[2][19][0] = 1'b1;
seq[2][19][1] = 1'b0;
seq[2][20][0] = 1'b0;
seq[2][20][1] = 1'b0;
seq[2][21][0] = 1'b1;
seq[2][21][1] = 1'b0;
seq[2][22][0] = 1'b1;
seq[2][22][1] = 1'b0;
seq[2][23][0] = 1'b1;
seq[2][23][1] = 1'b1;
seq[2][24][0] = 1'b0;
seq[2][24][1] = 1'b1;
seq[2][25][0] = 1'b0;
seq[2][25][1] = 1'b1;
seq[2][26][0] = 1'b1;
seq[2][26][1] = 1'b0;
seq[2][27][0] = 1'b1;
seq[2][27][1] = 1'b0;
seq[2][28][0] = 1'b1;
seq[2][28][1] = 1'b0;
seq[2][29][0] = 1'b1;
seq[2][29][1] = 1'b1;
seq[2][30][0] = 1'b0;
seq[2][30][1] = 1'b0;
seq[2][31][0] = 1'b0;
seq[2][31][1] = 1'b0;
seq[2][32][0] = 1'b0;
seq[2][32][1] = 1'b0;
seq[2][33][0] = 1'b0;
seq[2][33][1] = 1'b0;
seq[2][34][0] = 1'b1;
seq[2][34][1] = 1'b0;
seq[2][35][0] = 1'b1;
seq[2][35][1] = 1'b0;
seq[2][36][0] = 1'b1;
seq[2][36][1] = 1'b1;
seq[2][37][0] = 1'b1;
seq[2][37][1] = 1'b0;
seq[2][38][0] = 1'b1;
seq[2][38][1] = 1'b1;
seq[2][39][0] = 1'b1;
seq[2][39][1] = 1'b0;
seq[2][40][0] = 1'b0;
seq[2][40][1] = 1'b1;
seq[2][41][0] = 1'b0;
seq[2][41][1] = 1'b1;
seq[2][42][0] = 1'b1;
seq[2][42][1] = 1'b0;
seq[2][43][0] = 1'b0;
seq[2][43][1] = 1'b0;
seq[2][44][0] = 1'b0;
seq[2][44][1] = 1'b0;
seq[2][45][0] = 1'b1;
seq[2][45][1] = 1'b0;
seq[2][46][0] = 1'b1;
seq[2][46][1] = 1'b1;
seq[2][47][0] = 1'b1;
seq[2][47][1] = 1'b1;
seq[2][48][0] = 1'b1;
seq[2][48][1] = 1'b1;
seq[2][49][0] = 1'b1;
seq[2][49][1] = 1'b0;
seq[3][0][0] = 1'b0;
seq[3][0][1] = 1'b0;
seq[3][1][0] = 1'b0;
seq[3][1][1] = 1'b1;
seq[3][2][0] = 1'b0;
seq[3][2][1] = 1'b1;
seq[3][3][0] = 1'b0;
seq[3][3][1] = 1'b0;
seq[3][4][0] = 1'b1;
seq[3][4][1] = 1'b1;
seq[3][5][0] = 1'b1;
seq[3][5][1] = 1'b1;
seq[3][6][0] = 1'b0;
seq[3][6][1] = 1'b0;
seq[3][7][0] = 1'b0;
seq[3][7][1] = 1'b0;
seq[3][8][0] = 1'b1;
seq[3][8][1] = 1'b0;
seq[3][9][0] = 1'b1;
seq[3][9][1] = 1'b0;
seq[3][10][0] = 1'b1;
seq[3][10][1] = 1'b1;
seq[3][11][0] = 1'b0;
seq[3][11][1] = 1'b1;
seq[3][12][0] = 1'b1;
seq[3][12][1] = 1'b0;
seq[3][13][0] = 1'b0;
seq[3][13][1] = 1'b1;
seq[3][14][0] = 1'b1;
seq[3][14][1] = 1'b0;
seq[3][15][0] = 1'b0;
seq[3][15][1] = 1'b1;
seq[3][16][0] = 1'b0;
seq[3][16][1] = 1'b0;
seq[3][17][0] = 1'b1;
seq[3][17][1] = 1'b0;
seq[3][18][0] = 1'b1;
seq[3][18][1] = 1'b1;
seq[3][19][0] = 1'b0;
seq[3][19][1] = 1'b1;
seq[3][20][0] = 1'b0;
seq[3][20][1] = 1'b0;
seq[3][21][0] = 1'b1;
seq[3][21][1] = 1'b1;
seq[3][22][0] = 1'b0;
seq[3][22][1] = 1'b0;
seq[3][23][0] = 1'b0;
seq[3][23][1] = 1'b0;
seq[3][24][0] = 1'b0;
seq[3][24][1] = 1'b0;
seq[3][25][0] = 1'b1;
seq[3][25][1] = 1'b1;
seq[3][26][0] = 1'b0;
seq[3][26][1] = 1'b0;
seq[3][27][0] = 1'b0;
seq[3][27][1] = 1'b0;
seq[3][28][0] = 1'b0;
seq[3][28][1] = 1'b1;
seq[3][29][0] = 1'b0;
seq[3][29][1] = 1'b0;
seq[3][30][0] = 1'b1;
seq[3][30][1] = 1'b1;
seq[3][31][0] = 1'b0;
seq[3][31][1] = 1'b1;
seq[3][32][0] = 1'b1;
seq[3][32][1] = 1'b1;
seq[3][33][0] = 1'b0;
seq[3][33][1] = 1'b1;
seq[3][34][0] = 1'b0;
seq[3][34][1] = 1'b0;
seq[3][35][0] = 1'b1;
seq[3][35][1] = 1'b0;
seq[3][36][0] = 1'b0;
seq[3][36][1] = 1'b0;
seq[3][37][0] = 1'b1;
seq[3][37][1] = 1'b1;
seq[3][38][0] = 1'b0;
seq[3][38][1] = 1'b0;
seq[3][39][0] = 1'b0;
seq[3][39][1] = 1'b1;
seq[3][40][0] = 1'b0;
seq[3][40][1] = 1'b1;
seq[3][41][0] = 1'b1;
seq[3][41][1] = 1'b0;
seq[3][42][0] = 1'b1;
seq[3][42][1] = 1'b1;
seq[3][43][0] = 1'b1;
seq[3][43][1] = 1'b1;
seq[3][44][0] = 1'b1;
seq[3][44][1] = 1'b1;
seq[3][45][0] = 1'b0;
seq[3][45][1] = 1'b0;
seq[3][46][0] = 1'b1;
seq[3][46][1] = 1'b0;
seq[3][47][0] = 1'b1;
seq[3][47][1] = 1'b1;
seq[3][48][0] = 1'b1;
seq[3][48][1] = 1'b0;
seq[3][49][0] = 1'b1;
seq[3][49][1] = 1'b0;
seq[4][0][0] = 1'b0;
seq[4][0][1] = 1'b1;
seq[4][1][0] = 1'b1;
seq[4][1][1] = 1'b0;
seq[4][2][0] = 1'b1;
seq[4][2][1] = 1'b0;
seq[4][3][0] = 1'b1;
seq[4][3][1] = 1'b1;
seq[4][4][0] = 1'b0;
seq[4][4][1] = 1'b1;
seq[4][5][0] = 1'b0;
seq[4][5][1] = 1'b1;
seq[4][6][0] = 1'b1;
seq[4][6][1] = 1'b0;
seq[4][7][0] = 1'b0;
seq[4][7][1] = 1'b1;
seq[4][8][0] = 1'b0;
seq[4][8][1] = 1'b0;
seq[4][9][0] = 1'b1;
seq[4][9][1] = 1'b1;
seq[4][10][0] = 1'b0;
seq[4][10][1] = 1'b1;
seq[4][11][0] = 1'b1;
seq[4][11][1] = 1'b1;
seq[4][12][0] = 1'b1;
seq[4][12][1] = 1'b1;
seq[4][13][0] = 1'b1;
seq[4][13][1] = 1'b1;
seq[4][14][0] = 1'b1;
seq[4][14][1] = 1'b1;
seq[4][15][0] = 1'b0;
seq[4][15][1] = 1'b1;
seq[4][16][0] = 1'b1;
seq[4][16][1] = 1'b1;
seq[4][17][0] = 1'b1;
seq[4][17][1] = 1'b1;
seq[4][18][0] = 1'b1;
seq[4][18][1] = 1'b0;
seq[4][19][0] = 1'b1;
seq[4][19][1] = 1'b0;
seq[4][20][0] = 1'b1;
seq[4][20][1] = 1'b1;
seq[4][21][0] = 1'b1;
seq[4][21][1] = 1'b1;
seq[4][22][0] = 1'b1;
seq[4][22][1] = 1'b0;
seq[4][23][0] = 1'b1;
seq[4][23][1] = 1'b1;
seq[4][24][0] = 1'b0;
seq[4][24][1] = 1'b1;
seq[4][25][0] = 1'b0;
seq[4][25][1] = 1'b0;
seq[4][26][0] = 1'b0;
seq[4][26][1] = 1'b0;
seq[4][27][0] = 1'b1;
seq[4][27][1] = 1'b1;
seq[4][28][0] = 1'b1;
seq[4][28][1] = 1'b1;
seq[4][29][0] = 1'b1;
seq[4][29][1] = 1'b1;
seq[4][30][0] = 1'b1;
seq[4][30][1] = 1'b0;
seq[4][31][0] = 1'b1;
seq[4][31][1] = 1'b1;
seq[4][32][0] = 1'b0;
seq[4][32][1] = 1'b1;
seq[4][33][0] = 1'b0;
seq[4][33][1] = 1'b0;
seq[4][34][0] = 1'b1;
seq[4][34][1] = 1'b1;
seq[4][35][0] = 1'b0;
seq[4][35][1] = 1'b1;
seq[4][36][0] = 1'b1;
seq[4][36][1] = 1'b0;
seq[4][37][0] = 1'b1;
seq[4][37][1] = 1'b1;
seq[4][38][0] = 1'b1;
seq[4][38][1] = 1'b1;
seq[4][39][0] = 1'b0;
seq[4][39][1] = 1'b0;
seq[4][40][0] = 1'b0;
seq[4][40][1] = 1'b0;
seq[4][41][0] = 1'b1;
seq[4][41][1] = 1'b0;
seq[4][42][0] = 1'b1;
seq[4][42][1] = 1'b0;
seq[4][43][0] = 1'b1;
seq[4][43][1] = 1'b1;
seq[4][44][0] = 1'b1;
seq[4][44][1] = 1'b0;
seq[4][45][0] = 1'b0;
seq[4][45][1] = 1'b0;
seq[4][46][0] = 1'b1;
seq[4][46][1] = 1'b0;
seq[4][47][0] = 1'b0;
seq[4][47][1] = 1'b0;
seq[4][48][0] = 1'b0;
seq[4][48][1] = 1'b1;
seq[4][49][0] = 1'b1;
seq[4][49][1] = 1'b0;
seq[5][0][0] = 1'b1;
seq[5][0][1] = 1'b1;
seq[5][1][0] = 1'b0;
seq[5][1][1] = 1'b1;
seq[5][2][0] = 1'b1;
seq[5][2][1] = 1'b0;
seq[5][3][0] = 1'b0;
seq[5][3][1] = 1'b1;
seq[5][4][0] = 1'b1;
seq[5][4][1] = 1'b0;
seq[5][5][0] = 1'b0;
seq[5][5][1] = 1'b1;
seq[5][6][0] = 1'b1;
seq[5][6][1] = 1'b1;
seq[5][7][0] = 1'b0;
seq[5][7][1] = 1'b1;
seq[5][8][0] = 1'b1;
seq[5][8][1] = 1'b1;
seq[5][9][0] = 1'b1;
seq[5][9][1] = 1'b0;
seq[5][10][0] = 1'b1;
seq[5][10][1] = 1'b0;
seq[5][11][0] = 1'b1;
seq[5][11][1] = 1'b1;
seq[5][12][0] = 1'b0;
seq[5][12][1] = 1'b1;
seq[5][13][0] = 1'b1;
seq[5][13][1] = 1'b0;
seq[5][14][0] = 1'b1;
seq[5][14][1] = 1'b1;
seq[5][15][0] = 1'b0;
seq[5][15][1] = 1'b1;
seq[5][16][0] = 1'b0;
seq[5][16][1] = 1'b0;
seq[5][17][0] = 1'b0;
seq[5][17][1] = 1'b0;
seq[5][18][0] = 1'b0;
seq[5][18][1] = 1'b1;
seq[5][19][0] = 1'b1;
seq[5][19][1] = 1'b1;
seq[5][20][0] = 1'b1;
seq[5][20][1] = 1'b0;
seq[5][21][0] = 1'b1;
seq[5][21][1] = 1'b1;
seq[5][22][0] = 1'b0;
seq[5][22][1] = 1'b1;
seq[5][23][0] = 1'b1;
seq[5][23][1] = 1'b0;
seq[5][24][0] = 1'b1;
seq[5][24][1] = 1'b0;
seq[5][25][0] = 1'b0;
seq[5][25][1] = 1'b1;
seq[5][26][0] = 1'b1;
seq[5][26][1] = 1'b1;
seq[5][27][0] = 1'b1;
seq[5][27][1] = 1'b1;
seq[5][28][0] = 1'b1;
seq[5][28][1] = 1'b1;
seq[5][29][0] = 1'b0;
seq[5][29][1] = 1'b1;
seq[5][30][0] = 1'b1;
seq[5][30][1] = 1'b1;
seq[5][31][0] = 1'b0;
seq[5][31][1] = 1'b1;
seq[5][32][0] = 1'b0;
seq[5][32][1] = 1'b1;
seq[5][33][0] = 1'b0;
seq[5][33][1] = 1'b1;
seq[5][34][0] = 1'b0;
seq[5][34][1] = 1'b0;
seq[5][35][0] = 1'b1;
seq[5][35][1] = 1'b1;
seq[5][36][0] = 1'b0;
seq[5][36][1] = 1'b1;
seq[5][37][0] = 1'b0;
seq[5][37][1] = 1'b1;
seq[5][38][0] = 1'b1;
seq[5][38][1] = 1'b0;
seq[5][39][0] = 1'b0;
seq[5][39][1] = 1'b1;
seq[5][40][0] = 1'b1;
seq[5][40][1] = 1'b1;
seq[5][41][0] = 1'b1;
seq[5][41][1] = 1'b0;
seq[5][42][0] = 1'b1;
seq[5][42][1] = 1'b0;
seq[5][43][0] = 1'b1;
seq[5][43][1] = 1'b0;
seq[5][44][0] = 1'b1;
seq[5][44][1] = 1'b0;
seq[5][45][0] = 1'b0;
seq[5][45][1] = 1'b1;
seq[5][46][0] = 1'b0;
seq[5][46][1] = 1'b0;
seq[5][47][0] = 1'b0;
seq[5][47][1] = 1'b0;
seq[5][48][0] = 1'b1;
seq[5][48][1] = 1'b0;
seq[5][49][0] = 1'b1;
seq[5][49][1] = 1'b0;
seq[6][0][0] = 1'b1;
seq[6][0][1] = 1'b1;
seq[6][1][0] = 1'b0;
seq[6][1][1] = 1'b0;
seq[6][2][0] = 1'b1;
seq[6][2][1] = 1'b1;
seq[6][3][0] = 1'b0;
seq[6][3][1] = 1'b0;
seq[6][4][0] = 1'b0;
seq[6][4][1] = 1'b1;
seq[6][5][0] = 1'b0;
seq[6][5][1] = 1'b1;
seq[6][6][0] = 1'b0;
seq[6][6][1] = 1'b1;
seq[6][7][0] = 1'b1;
seq[6][7][1] = 1'b0;
seq[6][8][0] = 1'b0;
seq[6][8][1] = 1'b1;
seq[6][9][0] = 1'b1;
seq[6][9][1] = 1'b1;
seq[6][10][0] = 1'b0;
seq[6][10][1] = 1'b1;
seq[6][11][0] = 1'b0;
seq[6][11][1] = 1'b1;
seq[6][12][0] = 1'b0;
seq[6][12][1] = 1'b0;
seq[6][13][0] = 1'b0;
seq[6][13][1] = 1'b1;
seq[6][14][0] = 1'b1;
seq[6][14][1] = 1'b1;
seq[6][15][0] = 1'b0;
seq[6][15][1] = 1'b1;
seq[6][16][0] = 1'b1;
seq[6][16][1] = 1'b1;
seq[6][17][0] = 1'b0;
seq[6][17][1] = 1'b0;
seq[6][18][0] = 1'b1;
seq[6][18][1] = 1'b0;
seq[6][19][0] = 1'b1;
seq[6][19][1] = 1'b1;
seq[6][20][0] = 1'b1;
seq[6][20][1] = 1'b0;
seq[6][21][0] = 1'b0;
seq[6][21][1] = 1'b1;
seq[6][22][0] = 1'b1;
seq[6][22][1] = 1'b1;
seq[6][23][0] = 1'b1;
seq[6][23][1] = 1'b1;
seq[6][24][0] = 1'b1;
seq[6][24][1] = 1'b1;
seq[6][25][0] = 1'b0;
seq[6][25][1] = 1'b1;
seq[6][26][0] = 1'b1;
seq[6][26][1] = 1'b1;
seq[6][27][0] = 1'b1;
seq[6][27][1] = 1'b0;
seq[6][28][0] = 1'b0;
seq[6][28][1] = 1'b0;
seq[6][29][0] = 1'b0;
seq[6][29][1] = 1'b1;
seq[6][30][0] = 1'b1;
seq[6][30][1] = 1'b1;
seq[6][31][0] = 1'b0;
seq[6][31][1] = 1'b0;
seq[6][32][0] = 1'b0;
seq[6][32][1] = 1'b0;
seq[6][33][0] = 1'b0;
seq[6][33][1] = 1'b1;
seq[6][34][0] = 1'b1;
seq[6][34][1] = 1'b0;
seq[6][35][0] = 1'b0;
seq[6][35][1] = 1'b1;
seq[6][36][0] = 1'b0;
seq[6][36][1] = 1'b0;
seq[6][37][0] = 1'b0;
seq[6][37][1] = 1'b1;
seq[6][38][0] = 1'b1;
seq[6][38][1] = 1'b1;
seq[6][39][0] = 1'b1;
seq[6][39][1] = 1'b0;
seq[6][40][0] = 1'b1;
seq[6][40][1] = 1'b1;
seq[6][41][0] = 1'b1;
seq[6][41][1] = 1'b1;
seq[6][42][0] = 1'b1;
seq[6][42][1] = 1'b0;
seq[6][43][0] = 1'b1;
seq[6][43][1] = 1'b1;
seq[6][44][0] = 1'b0;
seq[6][44][1] = 1'b0;
seq[6][45][0] = 1'b0;
seq[6][45][1] = 1'b1;
seq[6][46][0] = 1'b1;
seq[6][46][1] = 1'b0;
seq[6][47][0] = 1'b0;
seq[6][47][1] = 1'b0;
seq[6][48][0] = 1'b0;
seq[6][48][1] = 1'b1;
seq[6][49][0] = 1'b1;
seq[6][49][1] = 1'b0;
seq[7][0][0] = 1'b1;
seq[7][0][1] = 1'b0;
seq[7][1][0] = 1'b1;
seq[7][1][1] = 1'b0;
seq[7][2][0] = 1'b1;
seq[7][2][1] = 1'b1;
seq[7][3][0] = 1'b0;
seq[7][3][1] = 1'b0;
seq[7][4][0] = 1'b0;
seq[7][4][1] = 1'b0;
seq[7][5][0] = 1'b0;
seq[7][5][1] = 1'b1;
seq[7][6][0] = 1'b0;
seq[7][6][1] = 1'b0;
seq[7][7][0] = 1'b1;
seq[7][7][1] = 1'b1;
seq[7][8][0] = 1'b1;
seq[7][8][1] = 1'b1;
seq[7][9][0] = 1'b1;
seq[7][9][1] = 1'b1;
seq[7][10][0] = 1'b1;
seq[7][10][1] = 1'b0;
seq[7][11][0] = 1'b1;
seq[7][11][1] = 1'b1;
seq[7][12][0] = 1'b0;
seq[7][12][1] = 1'b0;
seq[7][13][0] = 1'b0;
seq[7][13][1] = 1'b1;
seq[7][14][0] = 1'b0;
seq[7][14][1] = 1'b0;
seq[7][15][0] = 1'b0;
seq[7][15][1] = 1'b1;
seq[7][16][0] = 1'b1;
seq[7][16][1] = 1'b0;
seq[7][17][0] = 1'b1;
seq[7][17][1] = 1'b1;
seq[7][18][0] = 1'b0;
seq[7][18][1] = 1'b0;
seq[7][19][0] = 1'b1;
seq[7][19][1] = 1'b1;
seq[7][20][0] = 1'b1;
seq[7][20][1] = 1'b0;
seq[7][21][0] = 1'b1;
seq[7][21][1] = 1'b1;
seq[7][22][0] = 1'b0;
seq[7][22][1] = 1'b0;
seq[7][23][0] = 1'b0;
seq[7][23][1] = 1'b1;
seq[7][24][0] = 1'b0;
seq[7][24][1] = 1'b1;
seq[7][25][0] = 1'b0;
seq[7][25][1] = 1'b1;
seq[7][26][0] = 1'b1;
seq[7][26][1] = 1'b1;
seq[7][27][0] = 1'b1;
seq[7][27][1] = 1'b0;
seq[7][28][0] = 1'b0;
seq[7][28][1] = 1'b0;
seq[7][29][0] = 1'b1;
seq[7][29][1] = 1'b0;
seq[7][30][0] = 1'b1;
seq[7][30][1] = 1'b1;
seq[7][31][0] = 1'b0;
seq[7][31][1] = 1'b0;
seq[7][32][0] = 1'b0;
seq[7][32][1] = 1'b1;
seq[7][33][0] = 1'b1;
seq[7][33][1] = 1'b1;
seq[7][34][0] = 1'b0;
seq[7][34][1] = 1'b0;
seq[7][35][0] = 1'b0;
seq[7][35][1] = 1'b1;
seq[7][36][0] = 1'b1;
seq[7][36][1] = 1'b0;
seq[7][37][0] = 1'b0;
seq[7][37][1] = 1'b1;
seq[7][38][0] = 1'b1;
seq[7][38][1] = 1'b1;
seq[7][39][0] = 1'b1;
seq[7][39][1] = 1'b0;
seq[7][40][0] = 1'b0;
seq[7][40][1] = 1'b1;
seq[7][41][0] = 1'b1;
seq[7][41][1] = 1'b1;
seq[7][42][0] = 1'b1;
seq[7][42][1] = 1'b1;
seq[7][43][0] = 1'b0;
seq[7][43][1] = 1'b1;
seq[7][44][0] = 1'b1;
seq[7][44][1] = 1'b1;
seq[7][45][0] = 1'b1;
seq[7][45][1] = 1'b1;
seq[7][46][0] = 1'b0;
seq[7][46][1] = 1'b1;
seq[7][47][0] = 1'b1;
seq[7][47][1] = 1'b1;
seq[7][48][0] = 1'b1;
seq[7][48][1] = 1'b1;
seq[7][49][0] = 1'b0;
seq[7][49][1] = 1'b0;
seq[8][0][0] = 1'b1;
seq[8][0][1] = 1'b0;
seq[8][1][0] = 1'b0;
seq[8][1][1] = 1'b0;
seq[8][2][0] = 1'b1;
seq[8][2][1] = 1'b0;
seq[8][3][0] = 1'b1;
seq[8][3][1] = 1'b1;
seq[8][4][0] = 1'b1;
seq[8][4][1] = 1'b1;
seq[8][5][0] = 1'b0;
seq[8][5][1] = 1'b1;
seq[8][6][0] = 1'b1;
seq[8][6][1] = 1'b1;
seq[8][7][0] = 1'b1;
seq[8][7][1] = 1'b0;
seq[8][8][0] = 1'b1;
seq[8][8][1] = 1'b1;
seq[8][9][0] = 1'b1;
seq[8][9][1] = 1'b0;
seq[8][10][0] = 1'b1;
seq[8][10][1] = 1'b0;
seq[8][11][0] = 1'b1;
seq[8][11][1] = 1'b1;
seq[8][12][0] = 1'b1;
seq[8][12][1] = 1'b0;
seq[8][13][0] = 1'b1;
seq[8][13][1] = 1'b1;
seq[8][14][0] = 1'b0;
seq[8][14][1] = 1'b1;
seq[8][15][0] = 1'b0;
seq[8][15][1] = 1'b0;
seq[8][16][0] = 1'b0;
seq[8][16][1] = 1'b0;
seq[8][17][0] = 1'b1;
seq[8][17][1] = 1'b0;
seq[8][18][0] = 1'b0;
seq[8][18][1] = 1'b0;
seq[8][19][0] = 1'b0;
seq[8][19][1] = 1'b0;
seq[8][20][0] = 1'b1;
seq[8][20][1] = 1'b0;
seq[8][21][0] = 1'b1;
seq[8][21][1] = 1'b0;
seq[8][22][0] = 1'b1;
seq[8][22][1] = 1'b1;
seq[8][23][0] = 1'b0;
seq[8][23][1] = 1'b0;
seq[8][24][0] = 1'b1;
seq[8][24][1] = 1'b0;
seq[8][25][0] = 1'b1;
seq[8][25][1] = 1'b1;
seq[8][26][0] = 1'b1;
seq[8][26][1] = 1'b0;
seq[8][27][0] = 1'b0;
seq[8][27][1] = 1'b0;
seq[8][28][0] = 1'b1;
seq[8][28][1] = 1'b0;
seq[8][29][0] = 1'b1;
seq[8][29][1] = 1'b0;
seq[8][30][0] = 1'b0;
seq[8][30][1] = 1'b1;
seq[8][31][0] = 1'b1;
seq[8][31][1] = 1'b0;
seq[8][32][0] = 1'b1;
seq[8][32][1] = 1'b0;
seq[8][33][0] = 1'b0;
seq[8][33][1] = 1'b1;
seq[8][34][0] = 1'b0;
seq[8][34][1] = 1'b0;
seq[8][35][0] = 1'b1;
seq[8][35][1] = 1'b1;
seq[8][36][0] = 1'b0;
seq[8][36][1] = 1'b0;
seq[8][37][0] = 1'b1;
seq[8][37][1] = 1'b0;
seq[8][38][0] = 1'b1;
seq[8][38][1] = 1'b1;
seq[8][39][0] = 1'b0;
seq[8][39][1] = 1'b0;
seq[8][40][0] = 1'b1;
seq[8][40][1] = 1'b1;
seq[8][41][0] = 1'b1;
seq[8][41][1] = 1'b0;
seq[8][42][0] = 1'b1;
seq[8][42][1] = 1'b0;
seq[8][43][0] = 1'b0;
seq[8][43][1] = 1'b1;
seq[8][44][0] = 1'b1;
seq[8][44][1] = 1'b1;
seq[8][45][0] = 1'b0;
seq[8][45][1] = 1'b0;
seq[8][46][0] = 1'b1;
seq[8][46][1] = 1'b1;
seq[8][47][0] = 1'b1;
seq[8][47][1] = 1'b0;
seq[8][48][0] = 1'b1;
seq[8][48][1] = 1'b1;
seq[8][49][0] = 1'b1;
seq[8][49][1] = 1'b0;
seq[9][0][0] = 1'b1;
seq[9][0][1] = 1'b0;
seq[9][1][0] = 1'b0;
seq[9][1][1] = 1'b0;
seq[9][2][0] = 1'b1;
seq[9][2][1] = 1'b1;
seq[9][3][0] = 1'b1;
seq[9][3][1] = 1'b1;
seq[9][4][0] = 1'b1;
seq[9][4][1] = 1'b0;
seq[9][5][0] = 1'b0;
seq[9][5][1] = 1'b1;
seq[9][6][0] = 1'b0;
seq[9][6][1] = 1'b1;
seq[9][7][0] = 1'b0;
seq[9][7][1] = 1'b1;
seq[9][8][0] = 1'b1;
seq[9][8][1] = 1'b1;
seq[9][9][0] = 1'b1;
seq[9][9][1] = 1'b0;
seq[9][10][0] = 1'b1;
seq[9][10][1] = 1'b1;
seq[9][11][0] = 1'b1;
seq[9][11][1] = 1'b1;
seq[9][12][0] = 1'b1;
seq[9][12][1] = 1'b0;
seq[9][13][0] = 1'b1;
seq[9][13][1] = 1'b1;
seq[9][14][0] = 1'b1;
seq[9][14][1] = 1'b0;
seq[9][15][0] = 1'b0;
seq[9][15][1] = 1'b1;
seq[9][16][0] = 1'b1;
seq[9][16][1] = 1'b1;
seq[9][17][0] = 1'b0;
seq[9][17][1] = 1'b1;
seq[9][18][0] = 1'b1;
seq[9][18][1] = 1'b0;
seq[9][19][0] = 1'b1;
seq[9][19][1] = 1'b1;
seq[9][20][0] = 1'b0;
seq[9][20][1] = 1'b1;
seq[9][21][0] = 1'b1;
seq[9][21][1] = 1'b1;
seq[9][22][0] = 1'b1;
seq[9][22][1] = 1'b0;
seq[9][23][0] = 1'b0;
seq[9][23][1] = 1'b0;
seq[9][24][0] = 1'b1;
seq[9][24][1] = 1'b0;
seq[9][25][0] = 1'b1;
seq[9][25][1] = 1'b1;
seq[9][26][0] = 1'b0;
seq[9][26][1] = 1'b1;
seq[9][27][0] = 1'b0;
seq[9][27][1] = 1'b0;
seq[9][28][0] = 1'b0;
seq[9][28][1] = 1'b1;
seq[9][29][0] = 1'b0;
seq[9][29][1] = 1'b0;
seq[9][30][0] = 1'b0;
seq[9][30][1] = 1'b0;
seq[9][31][0] = 1'b0;
seq[9][31][1] = 1'b0;
seq[9][32][0] = 1'b1;
seq[9][32][1] = 1'b1;
seq[9][33][0] = 1'b1;
seq[9][33][1] = 1'b0;
seq[9][34][0] = 1'b1;
seq[9][34][1] = 1'b1;
seq[9][35][0] = 1'b1;
seq[9][35][1] = 1'b1;
seq[9][36][0] = 1'b1;
seq[9][36][1] = 1'b1;
seq[9][37][0] = 1'b0;
seq[9][37][1] = 1'b0;
seq[9][38][0] = 1'b1;
seq[9][38][1] = 1'b0;
seq[9][39][0] = 1'b1;
seq[9][39][1] = 1'b1;
seq[9][40][0] = 1'b1;
seq[9][40][1] = 1'b0;
seq[9][41][0] = 1'b1;
seq[9][41][1] = 1'b1;
seq[9][42][0] = 1'b1;
seq[9][42][1] = 1'b0;
seq[9][43][0] = 1'b0;
seq[9][43][1] = 1'b0;
seq[9][44][0] = 1'b0;
seq[9][44][1] = 1'b1;
seq[9][45][0] = 1'b0;
seq[9][45][1] = 1'b0;
seq[9][46][0] = 1'b1;
seq[9][46][1] = 1'b0;
seq[9][47][0] = 1'b0;
seq[9][47][1] = 1'b0;
seq[9][48][0] = 1'b1;
seq[9][48][1] = 1'b1;
seq[9][49][0] = 1'b1;
seq[9][49][1] = 1'b1;
seq[10][0][0] = 1'b0;
seq[10][0][1] = 1'b1;
seq[10][1][0] = 1'b1;
seq[10][1][1] = 1'b1;
seq[10][2][0] = 1'b1;
seq[10][2][1] = 1'b1;
seq[10][3][0] = 1'b1;
seq[10][3][1] = 1'b0;
seq[10][4][0] = 1'b0;
seq[10][4][1] = 1'b1;
seq[10][5][0] = 1'b0;
seq[10][5][1] = 1'b1;
seq[10][6][0] = 1'b1;
seq[10][6][1] = 1'b0;
seq[10][7][0] = 1'b0;
seq[10][7][1] = 1'b1;
seq[10][8][0] = 1'b1;
seq[10][8][1] = 1'b1;
seq[10][9][0] = 1'b1;
seq[10][9][1] = 1'b0;
seq[10][10][0] = 1'b1;
seq[10][10][1] = 1'b1;
seq[10][11][0] = 1'b0;
seq[10][11][1] = 1'b0;
seq[10][12][0] = 1'b1;
seq[10][12][1] = 1'b1;
seq[10][13][0] = 1'b0;
seq[10][13][1] = 1'b1;
seq[10][14][0] = 1'b0;
seq[10][14][1] = 1'b1;
seq[10][15][0] = 1'b1;
seq[10][15][1] = 1'b1;
seq[10][16][0] = 1'b1;
seq[10][16][1] = 1'b1;
seq[10][17][0] = 1'b1;
seq[10][17][1] = 1'b0;
seq[10][18][0] = 1'b1;
seq[10][18][1] = 1'b1;
seq[10][19][0] = 1'b0;
seq[10][19][1] = 1'b0;
seq[10][20][0] = 1'b0;
seq[10][20][1] = 1'b1;
seq[10][21][0] = 1'b0;
seq[10][21][1] = 1'b0;
seq[10][22][0] = 1'b1;
seq[10][22][1] = 1'b1;
seq[10][23][0] = 1'b0;
seq[10][23][1] = 1'b1;
seq[10][24][0] = 1'b0;
seq[10][24][1] = 1'b1;
seq[10][25][0] = 1'b1;
seq[10][25][1] = 1'b1;
seq[10][26][0] = 1'b0;
seq[10][26][1] = 1'b1;
seq[10][27][0] = 1'b0;
seq[10][27][1] = 1'b0;
seq[10][28][0] = 1'b0;
seq[10][28][1] = 1'b0;
seq[10][29][0] = 1'b0;
seq[10][29][1] = 1'b1;
seq[10][30][0] = 1'b0;
seq[10][30][1] = 1'b1;
seq[10][31][0] = 1'b0;
seq[10][31][1] = 1'b1;
seq[10][32][0] = 1'b0;
seq[10][32][1] = 1'b0;
seq[10][33][0] = 1'b1;
seq[10][33][1] = 1'b1;
seq[10][34][0] = 1'b1;
seq[10][34][1] = 1'b1;
seq[10][35][0] = 1'b1;
seq[10][35][1] = 1'b0;
seq[10][36][0] = 1'b0;
seq[10][36][1] = 1'b1;
seq[10][37][0] = 1'b0;
seq[10][37][1] = 1'b1;
seq[10][38][0] = 1'b0;
seq[10][38][1] = 1'b1;
seq[10][39][0] = 1'b1;
seq[10][39][1] = 1'b0;
seq[10][40][0] = 1'b0;
seq[10][40][1] = 1'b1;
seq[10][41][0] = 1'b0;
seq[10][41][1] = 1'b0;
seq[10][42][0] = 1'b0;
seq[10][42][1] = 1'b1;
seq[10][43][0] = 1'b1;
seq[10][43][1] = 1'b1;
seq[10][44][0] = 1'b1;
seq[10][44][1] = 1'b0;
seq[10][45][0] = 1'b1;
seq[10][45][1] = 1'b1;
seq[10][46][0] = 1'b0;
seq[10][46][1] = 1'b1;
seq[10][47][0] = 1'b1;
seq[10][47][1] = 1'b1;
seq[10][48][0] = 1'b1;
seq[10][48][1] = 1'b0;
seq[10][49][0] = 1'b0;
seq[10][49][1] = 1'b1;
seq[11][0][0] = 1'b1;
seq[11][0][1] = 1'b1;
seq[11][1][0] = 1'b1;
seq[11][1][1] = 1'b1;
seq[11][2][0] = 1'b0;
seq[11][2][1] = 1'b1;
seq[11][3][0] = 1'b1;
seq[11][3][1] = 1'b1;
seq[11][4][0] = 1'b0;
seq[11][4][1] = 1'b1;
seq[11][5][0] = 1'b0;
seq[11][5][1] = 1'b1;
seq[11][6][0] = 1'b0;
seq[11][6][1] = 1'b0;
seq[11][7][0] = 1'b1;
seq[11][7][1] = 1'b0;
seq[11][8][0] = 1'b1;
seq[11][8][1] = 1'b1;
seq[11][9][0] = 1'b1;
seq[11][9][1] = 1'b0;
seq[11][10][0] = 1'b0;
seq[11][10][1] = 1'b0;
seq[11][11][0] = 1'b1;
seq[11][11][1] = 1'b1;
seq[11][12][0] = 1'b1;
seq[11][12][1] = 1'b0;
seq[11][13][0] = 1'b1;
seq[11][13][1] = 1'b1;
seq[11][14][0] = 1'b1;
seq[11][14][1] = 1'b0;
seq[11][15][0] = 1'b1;
seq[11][15][1] = 1'b0;
seq[11][16][0] = 1'b0;
seq[11][16][1] = 1'b1;
seq[11][17][0] = 1'b0;
seq[11][17][1] = 1'b0;
seq[11][18][0] = 1'b0;
seq[11][18][1] = 1'b1;
seq[11][19][0] = 1'b0;
seq[11][19][1] = 1'b0;
seq[11][20][0] = 1'b1;
seq[11][20][1] = 1'b0;
seq[11][21][0] = 1'b1;
seq[11][21][1] = 1'b1;
seq[11][22][0] = 1'b1;
seq[11][22][1] = 1'b1;
seq[11][23][0] = 1'b0;
seq[11][23][1] = 1'b1;
seq[11][24][0] = 1'b0;
seq[11][24][1] = 1'b1;
seq[11][25][0] = 1'b1;
seq[11][25][1] = 1'b1;
seq[11][26][0] = 1'b0;
seq[11][26][1] = 1'b0;
seq[11][27][0] = 1'b0;
seq[11][27][1] = 1'b1;
seq[11][28][0] = 1'b0;
seq[11][28][1] = 1'b1;
seq[11][29][0] = 1'b1;
seq[11][29][1] = 1'b1;
seq[11][30][0] = 1'b0;
seq[11][30][1] = 1'b0;
seq[11][31][0] = 1'b0;
seq[11][31][1] = 1'b1;
seq[11][32][0] = 1'b0;
seq[11][32][1] = 1'b0;
seq[11][33][0] = 1'b0;
seq[11][33][1] = 1'b1;
seq[11][34][0] = 1'b1;
seq[11][34][1] = 1'b1;
seq[11][35][0] = 1'b1;
seq[11][35][1] = 1'b0;
seq[11][36][0] = 1'b0;
seq[11][36][1] = 1'b1;
seq[11][37][0] = 1'b0;
seq[11][37][1] = 1'b0;
seq[11][38][0] = 1'b1;
seq[11][38][1] = 1'b0;
seq[11][39][0] = 1'b1;
seq[11][39][1] = 1'b0;
seq[11][40][0] = 1'b0;
seq[11][40][1] = 1'b0;
seq[11][41][0] = 1'b1;
seq[11][41][1] = 1'b1;
seq[11][42][0] = 1'b0;
seq[11][42][1] = 1'b0;
seq[11][43][0] = 1'b1;
seq[11][43][1] = 1'b1;
seq[11][44][0] = 1'b1;
seq[11][44][1] = 1'b1;
seq[11][45][0] = 1'b1;
seq[11][45][1] = 1'b0;
seq[11][46][0] = 1'b1;
seq[11][46][1] = 1'b0;
seq[11][47][0] = 1'b0;
seq[11][47][1] = 1'b0;
seq[11][48][0] = 1'b0;
seq[11][48][1] = 1'b1;
seq[11][49][0] = 1'b1;
seq[11][49][1] = 1'b0;
seq[12][0][0] = 1'b1;
seq[12][0][1] = 1'b1;
seq[12][1][0] = 1'b1;
seq[12][1][1] = 1'b0;
seq[12][2][0] = 1'b0;
seq[12][2][1] = 1'b1;
seq[12][3][0] = 1'b1;
seq[12][3][1] = 1'b1;
seq[12][4][0] = 1'b1;
seq[12][4][1] = 1'b0;
seq[12][5][0] = 1'b0;
seq[12][5][1] = 1'b1;
seq[12][6][0] = 1'b0;
seq[12][6][1] = 1'b0;
seq[12][7][0] = 1'b0;
seq[12][7][1] = 1'b0;
seq[12][8][0] = 1'b1;
seq[12][8][1] = 1'b0;
seq[12][9][0] = 1'b0;
seq[12][9][1] = 1'b1;
seq[12][10][0] = 1'b1;
seq[12][10][1] = 1'b0;
seq[12][11][0] = 1'b0;
seq[12][11][1] = 1'b1;
seq[12][12][0] = 1'b0;
seq[12][12][1] = 1'b0;
seq[12][13][0] = 1'b1;
seq[12][13][1] = 1'b1;
seq[12][14][0] = 1'b1;
seq[12][14][1] = 1'b0;
seq[12][15][0] = 1'b0;
seq[12][15][1] = 1'b0;
seq[12][16][0] = 1'b0;
seq[12][16][1] = 1'b0;
seq[12][17][0] = 1'b0;
seq[12][17][1] = 1'b1;
seq[12][18][0] = 1'b0;
seq[12][18][1] = 1'b0;
seq[12][19][0] = 1'b1;
seq[12][19][1] = 1'b1;
seq[12][20][0] = 1'b0;
seq[12][20][1] = 1'b1;
seq[12][21][0] = 1'b0;
seq[12][21][1] = 1'b0;
seq[12][22][0] = 1'b1;
seq[12][22][1] = 1'b0;
seq[12][23][0] = 1'b1;
seq[12][23][1] = 1'b0;
seq[12][24][0] = 1'b0;
seq[12][24][1] = 1'b0;
seq[12][25][0] = 1'b0;
seq[12][25][1] = 1'b1;
seq[12][26][0] = 1'b0;
seq[12][26][1] = 1'b1;
seq[12][27][0] = 1'b0;
seq[12][27][1] = 1'b1;
seq[12][28][0] = 1'b0;
seq[12][28][1] = 1'b1;
seq[12][29][0] = 1'b1;
seq[12][29][1] = 1'b0;
seq[12][30][0] = 1'b1;
seq[12][30][1] = 1'b1;
seq[12][31][0] = 1'b1;
seq[12][31][1] = 1'b1;
seq[12][32][0] = 1'b1;
seq[12][32][1] = 1'b1;
seq[12][33][0] = 1'b0;
seq[12][33][1] = 1'b1;
seq[12][34][0] = 1'b0;
seq[12][34][1] = 1'b1;
seq[12][35][0] = 1'b0;
seq[12][35][1] = 1'b0;
seq[12][36][0] = 1'b1;
seq[12][36][1] = 1'b1;
seq[12][37][0] = 1'b1;
seq[12][37][1] = 1'b0;
seq[12][38][0] = 1'b0;
seq[12][38][1] = 1'b0;
seq[12][39][0] = 1'b0;
seq[12][39][1] = 1'b0;
seq[12][40][0] = 1'b1;
seq[12][40][1] = 1'b1;
seq[12][41][0] = 1'b0;
seq[12][41][1] = 1'b1;
seq[12][42][0] = 1'b0;
seq[12][42][1] = 1'b1;
seq[12][43][0] = 1'b1;
seq[12][43][1] = 1'b0;
seq[12][44][0] = 1'b0;
seq[12][44][1] = 1'b1;
seq[12][45][0] = 1'b1;
seq[12][45][1] = 1'b1;
seq[12][46][0] = 1'b1;
seq[12][46][1] = 1'b0;
seq[12][47][0] = 1'b1;
seq[12][47][1] = 1'b0;
seq[12][48][0] = 1'b0;
seq[12][48][1] = 1'b0;
seq[12][49][0] = 1'b0;
seq[12][49][1] = 1'b0;
seq[13][0][0] = 1'b1;
seq[13][0][1] = 1'b0;
seq[13][1][0] = 1'b1;
seq[13][1][1] = 1'b1;
seq[13][2][0] = 1'b1;
seq[13][2][1] = 1'b0;
seq[13][3][0] = 1'b0;
seq[13][3][1] = 1'b0;
seq[13][4][0] = 1'b0;
seq[13][4][1] = 1'b0;
seq[13][5][0] = 1'b1;
seq[13][5][1] = 1'b0;
seq[13][6][0] = 1'b1;
seq[13][6][1] = 1'b0;
seq[13][7][0] = 1'b0;
seq[13][7][1] = 1'b1;
seq[13][8][0] = 1'b0;
seq[13][8][1] = 1'b0;
seq[13][9][0] = 1'b1;
seq[13][9][1] = 1'b0;
seq[13][10][0] = 1'b0;
seq[13][10][1] = 1'b0;
seq[13][11][0] = 1'b0;
seq[13][11][1] = 1'b1;
seq[13][12][0] = 1'b1;
seq[13][12][1] = 1'b1;
seq[13][13][0] = 1'b0;
seq[13][13][1] = 1'b0;
seq[13][14][0] = 1'b0;
seq[13][14][1] = 1'b1;
seq[13][15][0] = 1'b0;
seq[13][15][1] = 1'b0;
seq[13][16][0] = 1'b1;
seq[13][16][1] = 1'b1;
seq[13][17][0] = 1'b1;
seq[13][17][1] = 1'b0;
seq[13][18][0] = 1'b1;
seq[13][18][1] = 1'b1;
seq[13][19][0] = 1'b1;
seq[13][19][1] = 1'b0;
seq[13][20][0] = 1'b1;
seq[13][20][1] = 1'b0;
seq[13][21][0] = 1'b0;
seq[13][21][1] = 1'b0;
seq[13][22][0] = 1'b1;
seq[13][22][1] = 1'b0;
seq[13][23][0] = 1'b1;
seq[13][23][1] = 1'b0;
seq[13][24][0] = 1'b0;
seq[13][24][1] = 1'b1;
seq[13][25][0] = 1'b0;
seq[13][25][1] = 1'b1;
seq[13][26][0] = 1'b0;
seq[13][26][1] = 1'b0;
seq[13][27][0] = 1'b0;
seq[13][27][1] = 1'b1;
seq[13][28][0] = 1'b1;
seq[13][28][1] = 1'b0;
seq[13][29][0] = 1'b0;
seq[13][29][1] = 1'b0;
seq[13][30][0] = 1'b0;
seq[13][30][1] = 1'b1;
seq[13][31][0] = 1'b1;
seq[13][31][1] = 1'b1;
seq[13][32][0] = 1'b1;
seq[13][32][1] = 1'b0;
seq[13][33][0] = 1'b0;
seq[13][33][1] = 1'b1;
seq[13][34][0] = 1'b1;
seq[13][34][1] = 1'b0;
seq[13][35][0] = 1'b1;
seq[13][35][1] = 1'b0;
seq[13][36][0] = 1'b1;
seq[13][36][1] = 1'b1;
seq[13][37][0] = 1'b0;
seq[13][37][1] = 1'b1;
seq[13][38][0] = 1'b1;
seq[13][38][1] = 1'b0;
seq[13][39][0] = 1'b0;
seq[13][39][1] = 1'b1;
seq[13][40][0] = 1'b0;
seq[13][40][1] = 1'b1;
seq[13][41][0] = 1'b0;
seq[13][41][1] = 1'b0;
seq[13][42][0] = 1'b1;
seq[13][42][1] = 1'b0;
seq[13][43][0] = 1'b0;
seq[13][43][1] = 1'b1;
seq[13][44][0] = 1'b1;
seq[13][44][1] = 1'b0;
seq[13][45][0] = 1'b0;
seq[13][45][1] = 1'b0;
seq[13][46][0] = 1'b0;
seq[13][46][1] = 1'b1;
seq[13][47][0] = 1'b1;
seq[13][47][1] = 1'b1;
seq[13][48][0] = 1'b1;
seq[13][48][1] = 1'b1;
seq[13][49][0] = 1'b1;
seq[13][49][1] = 1'b1;
seq[14][0][0] = 1'b0;
seq[14][0][1] = 1'b1;
seq[14][1][0] = 1'b0;
seq[14][1][1] = 1'b1;
seq[14][2][0] = 1'b1;
seq[14][2][1] = 1'b0;
seq[14][3][0] = 1'b0;
seq[14][3][1] = 1'b0;
seq[14][4][0] = 1'b0;
seq[14][4][1] = 1'b0;
seq[14][5][0] = 1'b1;
seq[14][5][1] = 1'b0;
seq[14][6][0] = 1'b0;
seq[14][6][1] = 1'b0;
seq[14][7][0] = 1'b0;
seq[14][7][1] = 1'b1;
seq[14][8][0] = 1'b0;
seq[14][8][1] = 1'b0;
seq[14][9][0] = 1'b1;
seq[14][9][1] = 1'b0;
seq[14][10][0] = 1'b1;
seq[14][10][1] = 1'b0;
seq[14][11][0] = 1'b1;
seq[14][11][1] = 1'b1;
seq[14][12][0] = 1'b1;
seq[14][12][1] = 1'b1;
seq[14][13][0] = 1'b1;
seq[14][13][1] = 1'b0;
seq[14][14][0] = 1'b0;
seq[14][14][1] = 1'b1;
seq[14][15][0] = 1'b1;
seq[14][15][1] = 1'b1;
seq[14][16][0] = 1'b0;
seq[14][16][1] = 1'b1;
seq[14][17][0] = 1'b1;
seq[14][17][1] = 1'b1;
seq[14][18][0] = 1'b0;
seq[14][18][1] = 1'b1;
seq[14][19][0] = 1'b0;
seq[14][19][1] = 1'b0;
seq[14][20][0] = 1'b0;
seq[14][20][1] = 1'b0;
seq[14][21][0] = 1'b1;
seq[14][21][1] = 1'b0;
seq[14][22][0] = 1'b1;
seq[14][22][1] = 1'b1;
seq[14][23][0] = 1'b0;
seq[14][23][1] = 1'b1;
seq[14][24][0] = 1'b1;
seq[14][24][1] = 1'b0;
seq[14][25][0] = 1'b0;
seq[14][25][1] = 1'b0;
seq[14][26][0] = 1'b0;
seq[14][26][1] = 1'b1;
seq[14][27][0] = 1'b1;
seq[14][27][1] = 1'b1;
seq[14][28][0] = 1'b1;
seq[14][28][1] = 1'b1;
seq[14][29][0] = 1'b1;
seq[14][29][1] = 1'b0;
seq[14][30][0] = 1'b0;
seq[14][30][1] = 1'b1;
seq[14][31][0] = 1'b1;
seq[14][31][1] = 1'b0;
seq[14][32][0] = 1'b1;
seq[14][32][1] = 1'b0;
seq[14][33][0] = 1'b1;
seq[14][33][1] = 1'b0;
seq[14][34][0] = 1'b1;
seq[14][34][1] = 1'b1;
seq[14][35][0] = 1'b1;
seq[14][35][1] = 1'b0;
seq[14][36][0] = 1'b0;
seq[14][36][1] = 1'b0;
seq[14][37][0] = 1'b0;
seq[14][37][1] = 1'b1;
seq[14][38][0] = 1'b1;
seq[14][38][1] = 1'b0;
seq[14][39][0] = 1'b0;
seq[14][39][1] = 1'b0;
seq[14][40][0] = 1'b1;
seq[14][40][1] = 1'b1;
seq[14][41][0] = 1'b1;
seq[14][41][1] = 1'b1;
seq[14][42][0] = 1'b1;
seq[14][42][1] = 1'b0;
seq[14][43][0] = 1'b1;
seq[14][43][1] = 1'b0;
seq[14][44][0] = 1'b1;
seq[14][44][1] = 1'b0;
seq[14][45][0] = 1'b0;
seq[14][45][1] = 1'b0;
seq[14][46][0] = 1'b1;
seq[14][46][1] = 1'b0;
seq[14][47][0] = 1'b1;
seq[14][47][1] = 1'b0;
seq[14][48][0] = 1'b1;
seq[14][48][1] = 1'b0;
seq[14][49][0] = 1'b0;
seq[14][49][1] = 1'b1;
seq[15][0][0] = 1'b1;
seq[15][0][1] = 1'b0;
seq[15][1][0] = 1'b1;
seq[15][1][1] = 1'b0;
seq[15][2][0] = 1'b0;
seq[15][2][1] = 1'b0;
seq[15][3][0] = 1'b0;
seq[15][3][1] = 1'b0;
seq[15][4][0] = 1'b1;
seq[15][4][1] = 1'b0;
seq[15][5][0] = 1'b0;
seq[15][5][1] = 1'b1;
seq[15][6][0] = 1'b0;
seq[15][6][1] = 1'b1;
seq[15][7][0] = 1'b0;
seq[15][7][1] = 1'b1;
seq[15][8][0] = 1'b0;
seq[15][8][1] = 1'b0;
seq[15][9][0] = 1'b1;
seq[15][9][1] = 1'b0;
seq[15][10][0] = 1'b0;
seq[15][10][1] = 1'b0;
seq[15][11][0] = 1'b1;
seq[15][11][1] = 1'b0;
seq[15][12][0] = 1'b0;
seq[15][12][1] = 1'b1;
seq[15][13][0] = 1'b0;
seq[15][13][1] = 1'b0;
seq[15][14][0] = 1'b0;
seq[15][14][1] = 1'b1;
seq[15][15][0] = 1'b1;
seq[15][15][1] = 1'b1;
seq[15][16][0] = 1'b1;
seq[15][16][1] = 1'b1;
seq[15][17][0] = 1'b1;
seq[15][17][1] = 1'b1;
seq[15][18][0] = 1'b1;
seq[15][18][1] = 1'b1;
seq[15][19][0] = 1'b0;
seq[15][19][1] = 1'b1;
seq[15][20][0] = 1'b1;
seq[15][20][1] = 1'b1;
seq[15][21][0] = 1'b0;
seq[15][21][1] = 1'b0;
seq[15][22][0] = 1'b1;
seq[15][22][1] = 1'b0;
seq[15][23][0] = 1'b1;
seq[15][23][1] = 1'b0;
seq[15][24][0] = 1'b0;
seq[15][24][1] = 1'b0;
seq[15][25][0] = 1'b0;
seq[15][25][1] = 1'b0;
seq[15][26][0] = 1'b0;
seq[15][26][1] = 1'b1;
seq[15][27][0] = 1'b1;
seq[15][27][1] = 1'b1;
seq[15][28][0] = 1'b1;
seq[15][28][1] = 1'b0;
seq[15][29][0] = 1'b0;
seq[15][29][1] = 1'b0;
seq[15][30][0] = 1'b0;
seq[15][30][1] = 1'b0;
seq[15][31][0] = 1'b1;
seq[15][31][1] = 1'b1;
seq[15][32][0] = 1'b1;
seq[15][32][1] = 1'b0;
seq[15][33][0] = 1'b0;
seq[15][33][1] = 1'b1;
seq[15][34][0] = 1'b1;
seq[15][34][1] = 1'b0;
seq[15][35][0] = 1'b1;
seq[15][35][1] = 1'b1;
seq[15][36][0] = 1'b0;
seq[15][36][1] = 1'b0;
seq[15][37][0] = 1'b0;
seq[15][37][1] = 1'b1;
seq[15][38][0] = 1'b1;
seq[15][38][1] = 1'b0;
seq[15][39][0] = 1'b1;
seq[15][39][1] = 1'b0;
seq[15][40][0] = 1'b1;
seq[15][40][1] = 1'b1;
seq[15][41][0] = 1'b0;
seq[15][41][1] = 1'b0;
seq[15][42][0] = 1'b0;
seq[15][42][1] = 1'b1;
seq[15][43][0] = 1'b1;
seq[15][43][1] = 1'b0;
seq[15][44][0] = 1'b0;
seq[15][44][1] = 1'b1;
seq[15][45][0] = 1'b1;
seq[15][45][1] = 1'b0;
seq[15][46][0] = 1'b1;
seq[15][46][1] = 1'b1;
seq[15][47][0] = 1'b0;
seq[15][47][1] = 1'b0;
seq[15][48][0] = 1'b1;
seq[15][48][1] = 1'b1;
seq[15][49][0] = 1'b0;
seq[15][49][1] = 1'b1;
seq[16][0][0] = 1'b1;
seq[16][0][1] = 1'b1;
seq[16][1][0] = 1'b1;
seq[16][1][1] = 1'b0;
seq[16][2][0] = 1'b0;
seq[16][2][1] = 1'b1;
seq[16][3][0] = 1'b0;
seq[16][3][1] = 1'b1;
seq[16][4][0] = 1'b0;
seq[16][4][1] = 1'b1;
seq[16][5][0] = 1'b1;
seq[16][5][1] = 1'b0;
seq[16][6][0] = 1'b0;
seq[16][6][1] = 1'b1;
seq[16][7][0] = 1'b0;
seq[16][7][1] = 1'b1;
seq[16][8][0] = 1'b1;
seq[16][8][1] = 1'b0;
seq[16][9][0] = 1'b0;
seq[16][9][1] = 1'b0;
seq[16][10][0] = 1'b1;
seq[16][10][1] = 1'b0;
seq[16][11][0] = 1'b0;
seq[16][11][1] = 1'b1;
seq[16][12][0] = 1'b1;
seq[16][12][1] = 1'b0;
seq[16][13][0] = 1'b1;
seq[16][13][1] = 1'b0;
seq[16][14][0] = 1'b1;
seq[16][14][1] = 1'b0;
seq[16][15][0] = 1'b1;
seq[16][15][1] = 1'b0;
seq[16][16][0] = 1'b0;
seq[16][16][1] = 1'b1;
seq[16][17][0] = 1'b1;
seq[16][17][1] = 1'b1;
seq[16][18][0] = 1'b1;
seq[16][18][1] = 1'b0;
seq[16][19][0] = 1'b1;
seq[16][19][1] = 1'b1;
seq[16][20][0] = 1'b1;
seq[16][20][1] = 1'b0;
seq[16][21][0] = 1'b1;
seq[16][21][1] = 1'b0;
seq[16][22][0] = 1'b1;
seq[16][22][1] = 1'b1;
seq[16][23][0] = 1'b0;
seq[16][23][1] = 1'b1;
seq[16][24][0] = 1'b1;
seq[16][24][1] = 1'b0;
seq[16][25][0] = 1'b1;
seq[16][25][1] = 1'b0;
seq[16][26][0] = 1'b1;
seq[16][26][1] = 1'b0;
seq[16][27][0] = 1'b1;
seq[16][27][1] = 1'b0;
seq[16][28][0] = 1'b1;
seq[16][28][1] = 1'b0;
seq[16][29][0] = 1'b0;
seq[16][29][1] = 1'b0;
seq[16][30][0] = 1'b0;
seq[16][30][1] = 1'b0;
seq[16][31][0] = 1'b0;
seq[16][31][1] = 1'b0;
seq[16][32][0] = 1'b1;
seq[16][32][1] = 1'b0;
seq[16][33][0] = 1'b1;
seq[16][33][1] = 1'b1;
seq[16][34][0] = 1'b1;
seq[16][34][1] = 1'b1;
seq[16][35][0] = 1'b0;
seq[16][35][1] = 1'b0;
seq[16][36][0] = 1'b1;
seq[16][36][1] = 1'b1;
seq[16][37][0] = 1'b0;
seq[16][37][1] = 1'b0;
seq[16][38][0] = 1'b0;
seq[16][38][1] = 1'b0;
seq[16][39][0] = 1'b0;
seq[16][39][1] = 1'b1;
seq[16][40][0] = 1'b0;
seq[16][40][1] = 1'b1;
seq[16][41][0] = 1'b1;
seq[16][41][1] = 1'b1;
seq[16][42][0] = 1'b1;
seq[16][42][1] = 1'b0;
seq[16][43][0] = 1'b1;
seq[16][43][1] = 1'b1;
seq[16][44][0] = 1'b1;
seq[16][44][1] = 1'b1;
seq[16][45][0] = 1'b0;
seq[16][45][1] = 1'b1;
seq[16][46][0] = 1'b0;
seq[16][46][1] = 1'b0;
seq[16][47][0] = 1'b0;
seq[16][47][1] = 1'b0;
seq[16][48][0] = 1'b0;
seq[16][48][1] = 1'b0;
seq[16][49][0] = 1'b0;
seq[16][49][1] = 1'b1;
seq[17][0][0] = 1'b1;
seq[17][0][1] = 1'b0;
seq[17][1][0] = 1'b0;
seq[17][1][1] = 1'b0;
seq[17][2][0] = 1'b1;
seq[17][2][1] = 1'b0;
seq[17][3][0] = 1'b0;
seq[17][3][1] = 1'b1;
seq[17][4][0] = 1'b0;
seq[17][4][1] = 1'b0;
seq[17][5][0] = 1'b1;
seq[17][5][1] = 1'b1;
seq[17][6][0] = 1'b1;
seq[17][6][1] = 1'b1;
seq[17][7][0] = 1'b1;
seq[17][7][1] = 1'b1;
seq[17][8][0] = 1'b1;
seq[17][8][1] = 1'b1;
seq[17][9][0] = 1'b1;
seq[17][9][1] = 1'b0;
seq[17][10][0] = 1'b0;
seq[17][10][1] = 1'b0;
seq[17][11][0] = 1'b1;
seq[17][11][1] = 1'b0;
seq[17][12][0] = 1'b1;
seq[17][12][1] = 1'b1;
seq[17][13][0] = 1'b1;
seq[17][13][1] = 1'b0;
seq[17][14][0] = 1'b1;
seq[17][14][1] = 1'b0;
seq[17][15][0] = 1'b0;
seq[17][15][1] = 1'b1;
seq[17][16][0] = 1'b0;
seq[17][16][1] = 1'b0;
seq[17][17][0] = 1'b1;
seq[17][17][1] = 1'b0;
seq[17][18][0] = 1'b0;
seq[17][18][1] = 1'b1;
seq[17][19][0] = 1'b1;
seq[17][19][1] = 1'b1;
seq[17][20][0] = 1'b0;
seq[17][20][1] = 1'b0;
seq[17][21][0] = 1'b0;
seq[17][21][1] = 1'b0;
seq[17][22][0] = 1'b1;
seq[17][22][1] = 1'b0;
seq[17][23][0] = 1'b0;
seq[17][23][1] = 1'b0;
seq[17][24][0] = 1'b1;
seq[17][24][1] = 1'b1;
seq[17][25][0] = 1'b0;
seq[17][25][1] = 1'b0;
seq[17][26][0] = 1'b1;
seq[17][26][1] = 1'b0;
seq[17][27][0] = 1'b0;
seq[17][27][1] = 1'b0;
seq[17][28][0] = 1'b1;
seq[17][28][1] = 1'b0;
seq[17][29][0] = 1'b1;
seq[17][29][1] = 1'b1;
seq[17][30][0] = 1'b0;
seq[17][30][1] = 1'b0;
seq[17][31][0] = 1'b0;
seq[17][31][1] = 1'b1;
seq[17][32][0] = 1'b0;
seq[17][32][1] = 1'b1;
seq[17][33][0] = 1'b1;
seq[17][33][1] = 1'b1;
seq[17][34][0] = 1'b0;
seq[17][34][1] = 1'b1;
seq[17][35][0] = 1'b0;
seq[17][35][1] = 1'b0;
seq[17][36][0] = 1'b0;
seq[17][36][1] = 1'b0;
seq[17][37][0] = 1'b0;
seq[17][37][1] = 1'b1;
seq[17][38][0] = 1'b0;
seq[17][38][1] = 1'b1;
seq[17][39][0] = 1'b1;
seq[17][39][1] = 1'b0;
seq[17][40][0] = 1'b1;
seq[17][40][1] = 1'b0;
seq[17][41][0] = 1'b1;
seq[17][41][1] = 1'b0;
seq[17][42][0] = 1'b0;
seq[17][42][1] = 1'b1;
seq[17][43][0] = 1'b0;
seq[17][43][1] = 1'b0;
seq[17][44][0] = 1'b1;
seq[17][44][1] = 1'b1;
seq[17][45][0] = 1'b1;
seq[17][45][1] = 1'b0;
seq[17][46][0] = 1'b0;
seq[17][46][1] = 1'b1;
seq[17][47][0] = 1'b1;
seq[17][47][1] = 1'b1;
seq[17][48][0] = 1'b0;
seq[17][48][1] = 1'b1;
seq[17][49][0] = 1'b1;
seq[17][49][1] = 1'b0;
seq[18][0][0] = 1'b1;
seq[18][0][1] = 1'b0;
seq[18][1][0] = 1'b1;
seq[18][1][1] = 1'b0;
seq[18][2][0] = 1'b1;
seq[18][2][1] = 1'b1;
seq[18][3][0] = 1'b1;
seq[18][3][1] = 1'b1;
seq[18][4][0] = 1'b0;
seq[18][4][1] = 1'b1;
seq[18][5][0] = 1'b0;
seq[18][5][1] = 1'b0;
seq[18][6][0] = 1'b0;
seq[18][6][1] = 1'b1;
seq[18][7][0] = 1'b0;
seq[18][7][1] = 1'b1;
seq[18][8][0] = 1'b1;
seq[18][8][1] = 1'b1;
seq[18][9][0] = 1'b0;
seq[18][9][1] = 1'b0;
seq[18][10][0] = 1'b1;
seq[18][10][1] = 1'b0;
seq[18][11][0] = 1'b1;
seq[18][11][1] = 1'b0;
seq[18][12][0] = 1'b0;
seq[18][12][1] = 1'b0;
seq[18][13][0] = 1'b0;
seq[18][13][1] = 1'b0;
seq[18][14][0] = 1'b0;
seq[18][14][1] = 1'b0;
seq[18][15][0] = 1'b0;
seq[18][15][1] = 1'b1;
seq[18][16][0] = 1'b0;
seq[18][16][1] = 1'b0;
seq[18][17][0] = 1'b1;
seq[18][17][1] = 1'b1;
seq[18][18][0] = 1'b0;
seq[18][18][1] = 1'b1;
seq[18][19][0] = 1'b0;
seq[18][19][1] = 1'b1;
seq[18][20][0] = 1'b1;
seq[18][20][1] = 1'b0;
seq[18][21][0] = 1'b1;
seq[18][21][1] = 1'b0;
seq[18][22][0] = 1'b0;
seq[18][22][1] = 1'b1;
seq[18][23][0] = 1'b1;
seq[18][23][1] = 1'b1;
seq[18][24][0] = 1'b1;
seq[18][24][1] = 1'b0;
seq[18][25][0] = 1'b0;
seq[18][25][1] = 1'b1;
seq[18][26][0] = 1'b0;
seq[18][26][1] = 1'b1;
seq[18][27][0] = 1'b0;
seq[18][27][1] = 1'b0;
seq[18][28][0] = 1'b0;
seq[18][28][1] = 1'b1;
seq[18][29][0] = 1'b0;
seq[18][29][1] = 1'b0;
seq[18][30][0] = 1'b0;
seq[18][30][1] = 1'b0;
seq[18][31][0] = 1'b1;
seq[18][31][1] = 1'b1;
seq[18][32][0] = 1'b0;
seq[18][32][1] = 1'b1;
seq[18][33][0] = 1'b1;
seq[18][33][1] = 1'b0;
seq[18][34][0] = 1'b1;
seq[18][34][1] = 1'b0;
seq[18][35][0] = 1'b1;
seq[18][35][1] = 1'b1;
seq[18][36][0] = 1'b1;
seq[18][36][1] = 1'b1;
seq[18][37][0] = 1'b0;
seq[18][37][1] = 1'b1;
seq[18][38][0] = 1'b1;
seq[18][38][1] = 1'b0;
seq[18][39][0] = 1'b0;
seq[18][39][1] = 1'b0;
seq[18][40][0] = 1'b1;
seq[18][40][1] = 1'b0;
seq[18][41][0] = 1'b1;
seq[18][41][1] = 1'b0;
seq[18][42][0] = 1'b1;
seq[18][42][1] = 1'b0;
seq[18][43][0] = 1'b0;
seq[18][43][1] = 1'b1;
seq[18][44][0] = 1'b1;
seq[18][44][1] = 1'b1;
seq[18][45][0] = 1'b1;
seq[18][45][1] = 1'b1;
seq[18][46][0] = 1'b0;
seq[18][46][1] = 1'b0;
seq[18][47][0] = 1'b0;
seq[18][47][1] = 1'b0;
seq[18][48][0] = 1'b0;
seq[18][48][1] = 1'b0;
seq[18][49][0] = 1'b1;
seq[18][49][1] = 1'b0;
seq[19][0][0] = 1'b1;
seq[19][0][1] = 1'b0;
seq[19][1][0] = 1'b1;
seq[19][1][1] = 1'b1;
seq[19][2][0] = 1'b0;
seq[19][2][1] = 1'b0;
seq[19][3][0] = 1'b1;
seq[19][3][1] = 1'b1;
seq[19][4][0] = 1'b1;
seq[19][4][1] = 1'b0;
seq[19][5][0] = 1'b0;
seq[19][5][1] = 1'b1;
seq[19][6][0] = 1'b0;
seq[19][6][1] = 1'b1;
seq[19][7][0] = 1'b1;
seq[19][7][1] = 1'b1;
seq[19][8][0] = 1'b1;
seq[19][8][1] = 1'b1;
seq[19][9][0] = 1'b1;
seq[19][9][1] = 1'b0;
seq[19][10][0] = 1'b1;
seq[19][10][1] = 1'b0;
seq[19][11][0] = 1'b1;
seq[19][11][1] = 1'b1;
seq[19][12][0] = 1'b1;
seq[19][12][1] = 1'b1;
seq[19][13][0] = 1'b1;
seq[19][13][1] = 1'b1;
seq[19][14][0] = 1'b1;
seq[19][14][1] = 1'b0;
seq[19][15][0] = 1'b0;
seq[19][15][1] = 1'b0;
seq[19][16][0] = 1'b1;
seq[19][16][1] = 1'b0;
seq[19][17][0] = 1'b0;
seq[19][17][1] = 1'b0;
seq[19][18][0] = 1'b0;
seq[19][18][1] = 1'b0;
seq[19][19][0] = 1'b1;
seq[19][19][1] = 1'b0;
seq[19][20][0] = 1'b1;
seq[19][20][1] = 1'b1;
seq[19][21][0] = 1'b0;
seq[19][21][1] = 1'b0;
seq[19][22][0] = 1'b0;
seq[19][22][1] = 1'b1;
seq[19][23][0] = 1'b1;
seq[19][23][1] = 1'b0;
seq[19][24][0] = 1'b1;
seq[19][24][1] = 1'b1;
seq[19][25][0] = 1'b1;
seq[19][25][1] = 1'b0;
seq[19][26][0] = 1'b1;
seq[19][26][1] = 1'b1;
seq[19][27][0] = 1'b1;
seq[19][27][1] = 1'b1;
seq[19][28][0] = 1'b1;
seq[19][28][1] = 1'b0;
seq[19][29][0] = 1'b0;
seq[19][29][1] = 1'b0;
seq[19][30][0] = 1'b1;
seq[19][30][1] = 1'b1;
seq[19][31][0] = 1'b0;
seq[19][31][1] = 1'b0;
seq[19][32][0] = 1'b0;
seq[19][32][1] = 1'b1;
seq[19][33][0] = 1'b0;
seq[19][33][1] = 1'b1;
seq[19][34][0] = 1'b0;
seq[19][34][1] = 1'b1;
seq[19][35][0] = 1'b0;
seq[19][35][1] = 1'b1;
seq[19][36][0] = 1'b0;
seq[19][36][1] = 1'b0;
seq[19][37][0] = 1'b1;
seq[19][37][1] = 1'b0;
seq[19][38][0] = 1'b1;
seq[19][38][1] = 1'b0;
seq[19][39][0] = 1'b1;
seq[19][39][1] = 1'b1;
seq[19][40][0] = 1'b0;
seq[19][40][1] = 1'b0;
seq[19][41][0] = 1'b0;
seq[19][41][1] = 1'b1;
seq[19][42][0] = 1'b1;
seq[19][42][1] = 1'b1;
seq[19][43][0] = 1'b1;
seq[19][43][1] = 1'b1;
seq[19][44][0] = 1'b1;
seq[19][44][1] = 1'b1;
seq[19][45][0] = 1'b1;
seq[19][45][1] = 1'b1;
seq[19][46][0] = 1'b0;
seq[19][46][1] = 1'b1;
seq[19][47][0] = 1'b1;
seq[19][47][1] = 1'b1;
seq[19][48][0] = 1'b1;
seq[19][48][1] = 1'b0;
seq[19][49][0] = 1'b1;
seq[19][49][1] = 1'b1;

end


endmodule